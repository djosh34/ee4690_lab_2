library ieee;

use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.math_real.all;

use std.textio.all;
use ieee.std_logic_textio.all;


package fc2_weights_package is
    constant HIDDEN_SIZE : integer := 608;
    constant OUTPUT_SIZE : integer := 10;

    type weights_2_type is array(0 to HIDDEN_SIZE - 1) of std_logic_vector(0 to OUTPUT_SIZE - 1);

    function read_and_populate_weights_2 return weights_2_type;
end fc2_weights_package;

package body fc2_weights_package is
    -- populate the weights_1 array
    function read_and_populate_weights_2 return weights_2_type is
      variable weights_array : weights_2_type;

    begin

      -- weights array: 608 x 10 
      -- weights_array(0) := "....";
      weights_array(0) := "1101010110";
      weights_array(1) := "0011000000";
      weights_array(2) := "0001110111";
      weights_array(3) := "0010110111";
      weights_array(4) := "1001100110";
      weights_array(5) := "0110101100";
      weights_array(6) := "1010111010";
      weights_array(7) := "1110100001";
      weights_array(8) := "1111100100";
      weights_array(9) := "0000111110";
      weights_array(10) := "1100101100";
      weights_array(11) := "1100111000";
      weights_array(12) := "1111000110";
      weights_array(13) := "0001110101";
      weights_array(14) := "1010000100";
      weights_array(15) := "1101100110";
      weights_array(16) := "1000110011";
      weights_array(17) := "0100001011";
      weights_array(18) := "1000010101";
      weights_array(19) := "1010011010";
      weights_array(20) := "0111100100";
      weights_array(21) := "1010000110";
      weights_array(22) := "0001110110";
      weights_array(23) := "1111110010";
      weights_array(24) := "0111001001";
      weights_array(25) := "1111000110";
      weights_array(26) := "0011010010";
      weights_array(27) := "0011111001";
      weights_array(28) := "1000101100";
      weights_array(29) := "0100111011";
      weights_array(30) := "1100101011";
      weights_array(31) := "1101011011";
      weights_array(32) := "0111000101";
      weights_array(33) := "1000101010";
      weights_array(34) := "1000001011";
      weights_array(35) := "0100000110";
      weights_array(36) := "1110010100";
      weights_array(37) := "1110101001";
      weights_array(38) := "0100110101";
      weights_array(39) := "0001011001";
      weights_array(40) := "1111000101";
      weights_array(41) := "0010010011";
      weights_array(42) := "1101010001";
      weights_array(43) := "0000110111";
      weights_array(44) := "1011010011";
      weights_array(45) := "0100101000";
      weights_array(46) := "1101101100";
      weights_array(47) := "0000111111";
      weights_array(48) := "1100011010";
      weights_array(49) := "1111000000";
      weights_array(50) := "1010110101";
      weights_array(51) := "1001111000";
      weights_array(52) := "1110010001";
      weights_array(53) := "0111000101";
      weights_array(54) := "1011100001";
      weights_array(55) := "0110011000";
      weights_array(56) := "1001110110";
      weights_array(57) := "1000101111";
      weights_array(58) := "1010011010";
      weights_array(59) := "1111000101";
      weights_array(60) := "0001110011";
      weights_array(61) := "1110110010";
      weights_array(62) := "1010100111";
      weights_array(63) := "0100101010";
      weights_array(64) := "1101101000";
      weights_array(65) := "0100101100";
      weights_array(66) := "1110001010";
      weights_array(67) := "1110011000";
      weights_array(68) := "1001011100";
      weights_array(69) := "0110011100";
      weights_array(70) := "1101110001";
      weights_array(71) := "1010010101";
      weights_array(72) := "0100001110";
      weights_array(73) := "1110100010";
      weights_array(74) := "1111011000";
      weights_array(75) := "0000011011";
      weights_array(76) := "0111011001";
      weights_array(77) := "1011000101";
      weights_array(78) := "1010101101";
      weights_array(79) := "0110000110";
      weights_array(80) := "1100001001";
      weights_array(81) := "1010001100";
      weights_array(82) := "0110100110";
      weights_array(83) := "0001100100";
      weights_array(84) := "0101101101";
      weights_array(85) := "0110101010";
      weights_array(86) := "0110010101";
      weights_array(87) := "0110101010";
      weights_array(88) := "0001001101";
      weights_array(89) := "0011100001";
      weights_array(90) := "1100101100";
      weights_array(91) := "1101010101";
      weights_array(92) := "1001001010";
      weights_array(93) := "1011110001";
      weights_array(94) := "1101101101";
      weights_array(95) := "0001111001";
      weights_array(96) := "1000011011";
      weights_array(97) := "0111000100";
      weights_array(98) := "0001001011";
      weights_array(99) := "0100011111";
      weights_array(100) := "0100111010";
      weights_array(101) := "1110000011";
      weights_array(102) := "1010101100";
      weights_array(103) := "1101100100";
      weights_array(104) := "1001100011";
      weights_array(105) := "0010101110";
      weights_array(106) := "0110011001";
      weights_array(107) := "1110000100";
      weights_array(108) := "1000011101";
      weights_array(109) := "0110011001";
      weights_array(110) := "0001111011";
      weights_array(111) := "0110101000";
      weights_array(112) := "0010000111";
      weights_array(113) := "0101010000";
      weights_array(114) := "0101101110";
      weights_array(115) := "1110101001";
      weights_array(116) := "1110000111";
      weights_array(117) := "1100001101";
      weights_array(118) := "0110100001";
      weights_array(119) := "0100011001";
      weights_array(120) := "0000111010";
      weights_array(121) := "1000001100";
      weights_array(122) := "0111100100";
      weights_array(123) := "0111011001";
      weights_array(124) := "0000101011";
      weights_array(125) := "1111001101";
      weights_array(126) := "0000011010";
      weights_array(127) := "0011001010";
      weights_array(128) := "0101110110";
      weights_array(129) := "1010001110";
      weights_array(130) := "0010101011";
      weights_array(131) := "0100001111";
      weights_array(132) := "0011011011";
      weights_array(133) := "0111000101";
      weights_array(134) := "1100100100";
      weights_array(135) := "0111111100";
      weights_array(136) := "1001001100";
      weights_array(137) := "1101101010";
      weights_array(138) := "0011011010";
      weights_array(139) := "1110100100";
      weights_array(140) := "0110000010";
      weights_array(141) := "1101011100";
      weights_array(142) := "1000111001";
      weights_array(143) := "1010111000";
      weights_array(144) := "1011010011";
      weights_array(145) := "0001011110";
      weights_array(146) := "1001011101";
      weights_array(147) := "1111010011";
      weights_array(148) := "1010010110";
      weights_array(149) := "1000010001";
      weights_array(150) := "0101100100";
      weights_array(151) := "0110100101";
      weights_array(152) := "0111001101";
      weights_array(153) := "1001101110";
      weights_array(154) := "0000110011";
      weights_array(155) := "0011001110";
      weights_array(156) := "0101111101";
      weights_array(157) := "1000101110";
      weights_array(158) := "1000100011";
      weights_array(159) := "0111101000";
      weights_array(160) := "1010111010";
      weights_array(161) := "0110011001";
      weights_array(162) := "0000111010";
      weights_array(163) := "1111000001";
      weights_array(164) := "1001000111";
      weights_array(165) := "0010101111";
      weights_array(166) := "0111001110";
      weights_array(167) := "1001100101";
      weights_array(168) := "1001001100";
      weights_array(169) := "0011010100";
      weights_array(170) := "1110010100";
      weights_array(171) := "1010111100";
      weights_array(172) := "1110011000";
      weights_array(173) := "0101100101";
      weights_array(174) := "0001110101";
      weights_array(175) := "0110001111";
      weights_array(176) := "0100100101";
      weights_array(177) := "0010100111";
      weights_array(178) := "1011100101";
      weights_array(179) := "1101000001";
      weights_array(180) := "0011100101";
      weights_array(181) := "0101111010";
      weights_array(182) := "1010100011";
      weights_array(183) := "0110000011";
      weights_array(184) := "1000111111";
      weights_array(185) := "0101000111";
      weights_array(186) := "1001101000";
      weights_array(187) := "0010010011";
      weights_array(188) := "0001110110";
      weights_array(189) := "0000110101";
      weights_array(190) := "0111101010";
      weights_array(191) := "1100101101";
      weights_array(192) := "0110001100";
      weights_array(193) := "1011101100";
      weights_array(194) := "0111000011";
      weights_array(195) := "0001011000";
      weights_array(196) := "0001110110";
      weights_array(197) := "1111011011";
      weights_array(198) := "1000010110";
      weights_array(199) := "0000111110";
      weights_array(200) := "1000101101";
      weights_array(201) := "1001010100";
      weights_array(202) := "1110101001";
      weights_array(203) := "1000111110";
      weights_array(204) := "1110100011";
      weights_array(205) := "1101100100";
      weights_array(206) := "0001110111";
      weights_array(207) := "1110101011";
      weights_array(208) := "1001000111";
      weights_array(209) := "0011101100";
      weights_array(210) := "0100100110";
      weights_array(211) := "1110110010";
      weights_array(212) := "0101111111";
      weights_array(213) := "1010000011";
      weights_array(214) := "0101010011";
      weights_array(215) := "0111000101";
      weights_array(216) := "0001011011";
      weights_array(217) := "0101011010";
      weights_array(218) := "0001111000";
      weights_array(219) := "1011011000";
      weights_array(220) := "1110100000";
      weights_array(221) := "1011001000";
      weights_array(222) := "1000100011";
      weights_array(223) := "1110000010";
      weights_array(224) := "1110001100";
      weights_array(225) := "0110010100";
      weights_array(226) := "0100001111";
      weights_array(227) := "1011001110";
      weights_array(228) := "1111000100";
      weights_array(229) := "1011100101";
      weights_array(230) := "0111001101";
      weights_array(231) := "0010110111";
      weights_array(232) := "1111100001";
      weights_array(233) := "1101001110";
      weights_array(234) := "1010110101";
      weights_array(235) := "1110101010";
      weights_array(236) := "1101000000";
      weights_array(237) := "0100000111";
      weights_array(238) := "0101011010";
      weights_array(239) := "0001010110";
      weights_array(240) := "0111100011";
      weights_array(241) := "0110001000";
      weights_array(242) := "0010101100";
      weights_array(243) := "0111011010";
      weights_array(244) := "1111011000";
      weights_array(245) := "0111100000";
      weights_array(246) := "0101100001";
      weights_array(247) := "1101011100";
      weights_array(248) := "0011100100";
      weights_array(249) := "1110010011";
      weights_array(250) := "1010101110";
      weights_array(251) := "1010110011";
      weights_array(252) := "0101101110";
      weights_array(253) := "0110010101";
      weights_array(254) := "1010001110";
      weights_array(255) := "1111101101";
      weights_array(256) := "1001100001";
      weights_array(257) := "0111000100";
      weights_array(258) := "1110011010";
      weights_array(259) := "0001110011";
      weights_array(260) := "0010110100";
      weights_array(261) := "0110111101";
      weights_array(262) := "0000110010";
      weights_array(263) := "0111011000";
      weights_array(264) := "0001110011";
      weights_array(265) := "0101110000";
      weights_array(266) := "1010100000";
      weights_array(267) := "1111000100";
      weights_array(268) := "1110000110";
      weights_array(269) := "0011010001";
      weights_array(270) := "1010001011";
      weights_array(271) := "1011000001";
      weights_array(272) := "0111101100";
      weights_array(273) := "0110100111";
      weights_array(274) := "0011001101";
      weights_array(275) := "1101100000";
      weights_array(276) := "1000111011";
      weights_array(277) := "0110010101";
      weights_array(278) := "0011110100";
      weights_array(279) := "0101110011";
      weights_array(280) := "1011000101";
      weights_array(281) := "0010111100";
      weights_array(282) := "0000011010";
      weights_array(283) := "1100101110";
      weights_array(284) := "1011110011";
      weights_array(285) := "1001011100";
      weights_array(286) := "1010011010";
      weights_array(287) := "0001101111";
      weights_array(288) := "0101100011";
      weights_array(289) := "1110011001";
      weights_array(290) := "1000000011";
      weights_array(291) := "1010111010";
      weights_array(292) := "0111010010";
      weights_array(293) := "1100101011";
      weights_array(294) := "0101001011";
      weights_array(295) := "0100100001";
      weights_array(296) := "1111001010";
      weights_array(297) := "0011111000";
      weights_array(298) := "0000111000";
      weights_array(299) := "1010101100";
      weights_array(300) := "1101011010";
      weights_array(301) := "0001100100";
      weights_array(302) := "1010011010";
      weights_array(303) := "0111111001";
      weights_array(304) := "0010100101";
      weights_array(305) := "0011000110";
      weights_array(306) := "0010101110";
      weights_array(307) := "0101110100";
      weights_array(308) := "0001011011";
      weights_array(309) := "1100101011";
      weights_array(310) := "0001010111";
      weights_array(311) := "1110001001";
      weights_array(312) := "1110001111";
      weights_array(313) := "0101010100";
      weights_array(314) := "1000101001";
      weights_array(315) := "1001101011";
      weights_array(316) := "1011110001";
      weights_array(317) := "1000111010";
      weights_array(318) := "1001111010";
      weights_array(319) := "1001100100";
      weights_array(320) := "1010011011";
      weights_array(321) := "0101111001";
      weights_array(322) := "0011010100";
      weights_array(323) := "1001010100";
      weights_array(324) := "0011101010";
      weights_array(325) := "1010110010";
      weights_array(326) := "1111000111";
      weights_array(327) := "0001111100";
      weights_array(328) := "0111011000";
      weights_array(329) := "0100110111";
      weights_array(330) := "0000000011";
      weights_array(331) := "0011001010";
      weights_array(332) := "1000111100";
      weights_array(333) := "1011110000";
      weights_array(334) := "1101011001";
      weights_array(335) := "0101010110";
      weights_array(336) := "1000100110";
      weights_array(337) := "1101111010";
      weights_array(338) := "1011101011";
      weights_array(339) := "1100011101";
      weights_array(340) := "0000010011";
      weights_array(341) := "1010111001";
      weights_array(342) := "0001000111";
      weights_array(343) := "0101001010";
      weights_array(344) := "0111101100";
      weights_array(345) := "1001101101";
      weights_array(346) := "0001001011";
      weights_array(347) := "0001111001";
      weights_array(348) := "0101000111";
      weights_array(349) := "1000011111";
      weights_array(350) := "1101110110";
      weights_array(351) := "0011011001";
      weights_array(352) := "1101001001";
      weights_array(353) := "0001110111";
      weights_array(354) := "0100111010";
      weights_array(355) := "1101111001";
      weights_array(356) := "1010001110";
      weights_array(357) := "1100010101";
      weights_array(358) := "1101000001";
      weights_array(359) := "1100110100";
      weights_array(360) := "1110001011";
      weights_array(361) := "1101010111";
      weights_array(362) := "0110101111";
      weights_array(363) := "0010111010";
      weights_array(364) := "1000101001";
      weights_array(365) := "0110101011";
      weights_array(366) := "1001011100";
      weights_array(367) := "1010001110";
      weights_array(368) := "0001010011";
      weights_array(369) := "0001001010";
      weights_array(370) := "0010011110";
      weights_array(371) := "0111010110";
      weights_array(372) := "0000101011";
      weights_array(373) := "0100111110";
      weights_array(374) := "1011010001";
      weights_array(375) := "1101100001";
      weights_array(376) := "0001110000";
      weights_array(377) := "0111001100";
      weights_array(378) := "0101011010";
      weights_array(379) := "1010001100";
      weights_array(380) := "1010101010";
      weights_array(381) := "1110111010";
      weights_array(382) := "0010110011";
      weights_array(383) := "1010001010";
      weights_array(384) := "1011001111";
      weights_array(385) := "1100011010";
      weights_array(386) := "1111010000";
      weights_array(387) := "0101000110";
      weights_array(388) := "0101101000";
      weights_array(389) := "0111011000";
      weights_array(390) := "0111101110";
      weights_array(391) := "1011100100";
      weights_array(392) := "1110101000";
      weights_array(393) := "1010011010";
      weights_array(394) := "0000111101";
      weights_array(395) := "0001001111";
      weights_array(396) := "1110100001";
      weights_array(397) := "0000111010";
      weights_array(398) := "0100100011";
      weights_array(399) := "0101111001";
      weights_array(400) := "0101010010";
      weights_array(401) := "1011010001";
      weights_array(402) := "0111111000";
      weights_array(403) := "1110101110";
      weights_array(404) := "0110110001";
      weights_array(405) := "0110001100";
      weights_array(406) := "1111100000";
      weights_array(407) := "0011100010";
      weights_array(408) := "0011100011";
      weights_array(409) := "1011110100";
      weights_array(410) := "0110110011";
      weights_array(411) := "1100000101";
      weights_array(412) := "0000110001";
      weights_array(413) := "0110110010";
      weights_array(414) := "0111100010";
      weights_array(415) := "1110110001";
      weights_array(416) := "0010111111";
      weights_array(417) := "1010010010";
      weights_array(418) := "1100100010";
      weights_array(419) := "1001001010";
      weights_array(420) := "1101001001";
      weights_array(421) := "0011010011";
      weights_array(422) := "1001001110";
      weights_array(423) := "0111001100";
      weights_array(424) := "1010100110";
      weights_array(425) := "1010100011";
      weights_array(426) := "0011110101";
      weights_array(427) := "1111111011";
      weights_array(428) := "0011110011";
      weights_array(429) := "0111100010";
      weights_array(430) := "0111011110";
      weights_array(431) := "1101001011";
      weights_array(432) := "0100010101";
      weights_array(433) := "0010100101";
      weights_array(434) := "0111110010";
      weights_array(435) := "0101111100";
      weights_array(436) := "1101011001";
      weights_array(437) := "1010110001";
      weights_array(438) := "1011011010";
      weights_array(439) := "0111000100";
      weights_array(440) := "1000100101";
      weights_array(441) := "0110001110";
      weights_array(442) := "0000010110";
      weights_array(443) := "0010100011";
      weights_array(444) := "0101101000";
      weights_array(445) := "0010111100";
      weights_array(446) := "0011001101";
      weights_array(447) := "0101110101";
      weights_array(448) := "0011010010";
      weights_array(449) := "0110000001";
      weights_array(450) := "0100011011";
      weights_array(451) := "1000110011";
      weights_array(452) := "0110001000";
      weights_array(453) := "1001001101";
      weights_array(454) := "0001010111";
      weights_array(455) := "1101110001";
      weights_array(456) := "1100011001";
      weights_array(457) := "1010100011";
      weights_array(458) := "0101000110";
      weights_array(459) := "1111110100";
      weights_array(460) := "1100010110";
      weights_array(461) := "1101010101";
      weights_array(462) := "1011000100";
      weights_array(463) := "0101010010";
      weights_array(464) := "1111001010";
      weights_array(465) := "1000001101";
      weights_array(466) := "0010101110";
      weights_array(467) := "0101000110";
      weights_array(468) := "1001001011";
      weights_array(469) := "1111001101";
      weights_array(470) := "0011100110";
      weights_array(471) := "1101011111";
      weights_array(472) := "0100000111";
      weights_array(473) := "1011111000";
      weights_array(474) := "0011000110";
      weights_array(475) := "1111001111";
      weights_array(476) := "1100001101";
      weights_array(477) := "1001001111";
      weights_array(478) := "0101101001";
      weights_array(479) := "1111101000";
      weights_array(480) := "0000111001";
      weights_array(481) := "0000011110";
      weights_array(482) := "1000010011";
      weights_array(483) := "0000101011";
      weights_array(484) := "0100111011";
      weights_array(485) := "0111001000";
      weights_array(486) := "1010010101";
      weights_array(487) := "1000001001";
      weights_array(488) := "1001011000";
      weights_array(489) := "1111110010";
      weights_array(490) := "0010011101";
      weights_array(491) := "0010101001";
      weights_array(492) := "0011100111";
      weights_array(493) := "1110100000";
      weights_array(494) := "1000100011";
      weights_array(495) := "1000111100";
      weights_array(496) := "0101010001";
      weights_array(497) := "1100101011";
      weights_array(498) := "0111000011";
      weights_array(499) := "0001110101";
      weights_array(500) := "0000111100";
      weights_array(501) := "0001011101";
      weights_array(502) := "1001011010";
      weights_array(503) := "0111100100";
      weights_array(504) := "1110100110";
      weights_array(505) := "0111001000";
      weights_array(506) := "0110110100";
      weights_array(507) := "1101101000";
      weights_array(508) := "0100010111";
      weights_array(509) := "1011011101";
      weights_array(510) := "1100010100";
      weights_array(511) := "0111010011";
      weights_array(512) := "1011110110";
      weights_array(513) := "1010010110";
      weights_array(514) := "1101111010";
      weights_array(515) := "1000100001";
      weights_array(516) := "1011010100";
      weights_array(517) := "1101001101";
      weights_array(518) := "1111000001";
      weights_array(519) := "1010001101";
      weights_array(520) := "0010011000";
      weights_array(521) := "1011010110";
      weights_array(522) := "1000100110";
      weights_array(523) := "0111110100";
      weights_array(524) := "0110000011";
      weights_array(525) := "0110011000";
      weights_array(526) := "1010001001";
      weights_array(527) := "0101010110";
      weights_array(528) := "1110111010";
      weights_array(529) := "1101111100";
      weights_array(530) := "0111100010";
      weights_array(531) := "0111100111";
      weights_array(532) := "1000011110";
      weights_array(533) := "0000101111";
      weights_array(534) := "0110100010";
      weights_array(535) := "0110010010";
      weights_array(536) := "1111100110";
      weights_array(537) := "0010100010";
      weights_array(538) := "1000111010";
      weights_array(539) := "1001011101";
      weights_array(540) := "1011001100";
      weights_array(541) := "1111001000";
      weights_array(542) := "0011010110";
      weights_array(543) := "0101010010";
      weights_array(544) := "1110001100";
      weights_array(545) := "0010000011";
      weights_array(546) := "1101010110";
      weights_array(547) := "1000101111";
      weights_array(548) := "1000101001";
      weights_array(549) := "0100101100";
      weights_array(550) := "1110001000";
      weights_array(551) := "1111011100";
      weights_array(552) := "0001101011";
      weights_array(553) := "0101010001";
      weights_array(554) := "1000011010";
      weights_array(555) := "1101100010";
      weights_array(556) := "0111010001";
      weights_array(557) := "1100111100";
      weights_array(558) := "1101011001";
      weights_array(559) := "0111101001";
      weights_array(560) := "1001101101";
      weights_array(561) := "1011001111";
      weights_array(562) := "0010011100";
      weights_array(563) := "0100110100";
      weights_array(564) := "1101000010";
      weights_array(565) := "0110100111";
      weights_array(566) := "1100110100";
      weights_array(567) := "1101111000";
      weights_array(568) := "0100011010";
      weights_array(569) := "1011100111";
      weights_array(570) := "1010110101";
      weights_array(571) := "0011100100";
      weights_array(572) := "1111000100";
      weights_array(573) := "0111110100";
      weights_array(574) := "1010100110";
      weights_array(575) := "0110010001";
      weights_array(576) := "1100000111";
      weights_array(577) := "1110001100";
      weights_array(578) := "1000011011";
      weights_array(579) := "0011100111";
      weights_array(580) := "0010000001";
      weights_array(581) := "0111110100";
      weights_array(582) := "1110111110";
      weights_array(583) := "1000100001";
      weights_array(584) := "0101011100";
      weights_array(585) := "0100100100";
      weights_array(586) := "0000101101";
      weights_array(587) := "0110101011";
      weights_array(588) := "1001000101";
      weights_array(589) := "0100110011";
      weights_array(590) := "1110101010";
      weights_array(591) := "0010010011";
      weights_array(592) := "1001000101";
      weights_array(593) := "0100011011";
      weights_array(594) := "0111100101";
      weights_array(595) := "0101100100";
      weights_array(596) := "1011100101";
      weights_array(597) := "1001101101";
      weights_array(598) := "1000011100";
      weights_array(599) := "0110000100";
      weights_array(600) := "0000001101";
      weights_array(601) := "0011110000";
      weights_array(602) := "0001100010";
      weights_array(603) := "0011111100";
      weights_array(604) := "0011011100";
      weights_array(605) := "1010110110";
      weights_array(606) := "1100111010";
      weights_array(607) := "1001100001";

      return weights_array;
    end function;
end fc2_weights_package;

