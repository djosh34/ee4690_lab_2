library ieee;

use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.math_real.all;

use std.textio.all;
use ieee.std_logic_textio.all;


package fc2_weights_package is
    constant HIDDEN_SIZE : integer := 608;
    constant OUTPUT_SIZE : integer := 10;

    type weights_2_type is array(0 to HIDDEN_SIZE - 1) of std_logic_vector(0 to OUTPUT_SIZE - 1);

    function read_and_populate_weights_2 return weights_2_type;
end fc2_weights_package;

package body fc2_weights_package is
    -- populate the weights_1 array
    function read_and_populate_weights_2 return weights_2_type is
      variable weights_array : weights_2_type;

    begin

      -- weights array: 608 x 768 
      -- weights_array(0) := "....";
            weights_array(0) := "10001011101110111011010101001011011011001010101011111010111101101011101101100110110000000011111010000111100110000001110001000100010000101101011110111100010001101001100110111000001100101010000101000110111111011001010000011111100111001111100000001001011100111010000000111011000110001001111001110100100110100000010110111111100101100000111011110100010001101001111111001011000000110001110111100001110010000101001001010001011110101101000100001110100000000001010111011110110011010101110100100011110001110100001010010110111111110110001011001000101111001011101100110110110010110110101011100011000010101000111000000111";
      weights_array(1) := "10000101101110010100100111000111100111101010011011001101000101011111011011101001101011110011001001011101001101010111111100110100100101110101110000010011100010010101001000101101100101010100001110100100001011010011101101001001111010101101111011011111010011010110010101011000110101010001000011001111100010010001010111000000010000101100001101010001100010101011011111100100000101010110010001111110100010111011111000110111001010010001011110111001010010010110100110111101100101011001101100001100010001001110000111111011001001100001110111110011100001011010011101011111000111111000110111000110110101100111000100000010";
      weights_array(2) := "01010111100010100001110111110000100011001100100001101111001101100011010101101111011001110100010001000110011101011001101000110101011011010011100110011001100100011101011001111001011010110001001011100100001010010101010100011101110111111011000011111100111101110110110100111111111001101100101001011000110100111110000110001000101011101001010000100100100000010000100010110101001100100101111110100111110010000111111111100111110001011111111001100111010101101100100001010010101001100111000100000110011111000010000111100101110010111101111010110011110011101100001100001001011001000111111101011110000100110010100101011100";
      weights_array(3) := "11101000100011010000101111110001100000011010101001010110100110001000101000101100000110001101111101100001100000100110000000110101100011011110010011110010110110010001101111000110001111000110101001111100010001101100101111110100000111101100101110011111100010011101000111010101101100111000110110001010110011010101101001011011011110111001011101100011111110111101001001000010110100111110000010111111000100011110001111000010000111110011111100111011000010111000011100110111100111110111011100000100110010001011011101010101101011100101000101110000100111110010000111011011110010010101110000010100100010001011110001111001";
      weights_array(4) := "00111111111101011000101100011110010001100001011100110010110011111100001001000010001111010110011100001011110000110011001010101000101000110101001100000011011011111010010100010110111011101010111101001001101111110111100000101010000001011011000010100110101110011001111011100000110110110101100110010101011101011011010000111111010011010100110011100100110100100111000100111100000011011000111000001011101011110011101111101111101000001111110001110100100111010001000101010000001000100100001110011000010111110101100110110000101100000011000011110110111000000001110010010101100101110111011000010111011101100011110001110111";
      weights_array(5) := "10110010010101001011001100110101000010110111100110111001101011000001111100111000000000100001010110011000001011100100000110010010100010010010011111111100001010001110000001111010000001001001110000011111010100100001101011110000010000010010001100011001010101000011111111000100000011110110111001011000011010110001101001001110111101011100111101011100000101110111010101010010101101101010011001100100011001011110100001101101110001000011101010111110001001011011001110011101000000010100000011101010111000011001111000101111111010001101010111001001001100110010000101101110001100111010010100100110100001010100001001011110";
      weights_array(6) := "00000110011100000101000010011111011001010000011110010001011000011111110010111010110011011010101110111010011011110011010111011111011110011110011101100000110111011110011010011001000001001010001111010101101100010100100011110100101100100101001001111001001010110010010100000010101010000111011101010110111110110010110110110110110010011001101001110101111101011011100010111111011011000111110111001110111101010011010000000000100110110001001100011010010011100010110010000000111011010101111111011101101100010100111001010100001001011000011011001100001111001001111110100111111000011000000001100010101100100100011010011010";
      weights_array(7) := "10111100111011110010111001001000100110101001001100100100110100100100110110000111011110101011001001010011010110001010110001100100110101111001010001101011110111000000111111110111111010001100110111001011110101101110100100000000111111110110010100100001101011110100110000011000111001101101010100000000000101001111001011000001001100110100100110010010110011100100110101100011001101000101000010010011001100000001010001010000100000111010001011010001111001110000011000111110011101111011110001000010001010010001110110101110110011010111000101011100100110101011010100000100111101100111111011010110111010001011111110011100";
      weights_array(8) := "10111010010010011101011101100111011100000101100110000000111011110010000011010001001001010000100010111100110000101010100010001011111110000110100011011000011101101010111000000001010001111101101000101111000110111011111011000011001100010101011110010000011110100011001010001010010010010011101110111110100010100110111010010110100011100111000111101011001011100110100011110101111111000010111111010010010101101001000110100110111101101101111100100010011100001011001001101001101110111011010001111000010010100110001010001001111000000110100110111111111000110111000010110000010011001100001010110010000101110100000000100110";
      weights_array(9) := "00110001000001001110000010010111101001111111100100101110010110100000001100011110100010101101011110110100101011101001111100011100001111000000001010110101101010100101110100000111111110111101010100100100101010111000111110000010001001111010010010000010010101011001010010000111011011011000100111100111000000011000111110111000110000100110001000111110011111011101011011101100100010110000001010000000001110110100100010111001100011000111100111001100100100110111011111000100010011011001111010111011001110101111010000001101000101110000101000010100000100000101100011001011110001000110000110111001001111011110110010000001";

      return weights_array;
    end function;
end fc2_weights_package;

