library ieee;

use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.math_real.all;

use std.textio.all;
use ieee.std_logic_textio.all;


package fc2_weights_package is
    constant HIDDEN_SIZE : integer := 608;
    constant OUTPUT_SIZE : integer := 10;

    type weights_2_type is array(0 to HIDDEN_SIZE - 1) of std_logic_vector(0 to OUTPUT_SIZE - 1);

    function read_and_populate_weights_2 return weights_2_type;
end fc2_weights_package;

package body fc2_weights_package is
    -- populate the weights_1 array
    function read_and_populate_weights_2 return weights_2_type is
      variable weights_array : weights_2_type;

    begin

      -- weights array: 608 x 768 
      -- weights_array(0) := "....";
      weights_array(0) := "1110101000";
      weights_array(1) := "1101000110";
      weights_array(2) := "0001010001";
      weights_array(3) := "0100000111";
      weights_array(4) := "0101100001";
      weights_array(5) := "1110001100";
      weights_array(6) := "1011000001";
      weights_array(7) := "1011010000";
      weights_array(8) := "0100001101";
      weights_array(9) := "1011010001";
      weights_array(10) := "1100001101";
      weights_array(11) := "0110100111";
      weights_array(12) := "0011110011";
      weights_array(13) := "0110100111";
      weights_array(14) := "1010001100";
      weights_array(15) := "0111101000";
      weights_array(16) := "1010010010";
      weights_array(17) := "1000101100";
      weights_array(18) := "1100011101";
      weights_array(19) := "0111010010";
      weights_array(20) := "0110101010";
      weights_array(21) := "1010010110";
      weights_array(22) := "0100101110";
      weights_array(23) := "1000101100";
      weights_array(24) := "1101010100";
      weights_array(25) := "0110010001";
      weights_array(26) := "0111000110";
      weights_array(27) := "1001011000";
      weights_array(28) := "1100011110";
      weights_array(29) := "0101110100";
      weights_array(30) := "0100100101";
      weights_array(31) := "0111101000";
      weights_array(32) := "0101100010";
      weights_array(33) := "0000010001";
      weights_array(34) := "0001110001";
      weights_array(35) := "0011010100";
      weights_array(36) := "0011101010";
      weights_array(37) := "1001011100";
      weights_array(38) := "0110100011";
      weights_array(39) := "1101010100";
      weights_array(40) := "0111000010";
      weights_array(41) := "1010001110";
      weights_array(42) := "0111110000";
      weights_array(43) := "0011101101";
      weights_array(44) := "0011010110";
      weights_array(45) := "0001000100";
      weights_array(46) := "1011010001";
      weights_array(47) := "0011010010";
      weights_array(48) := "1111001000";
      weights_array(49) := "1010011110";
      weights_array(50) := "0011100110";
      weights_array(51) := "0101010010";
      weights_array(52) := "1011010100";
      weights_array(53) := "0010101100";
      weights_array(54) := "0001111110";
      weights_array(55) := "1011010101";
      weights_array(56) := "0010010110";
      weights_array(57) := "1011001001";
      weights_array(58) := "0101100101";
      weights_array(59) := "1010100100";
      weights_array(60) := "0011001001";
      weights_array(61) := "1101100100";
      weights_array(62) := "1010101000";
      weights_array(63) := "1011101000";
      weights_array(64) := "1010111010";
      weights_array(65) := "1000011111";
      weights_array(66) := "1000110111";
      weights_array(67) := "0011001111";
      weights_array(68) := "1001000101";
      weights_array(69) := "0001111101";
      weights_array(70) := "1011000101";
      weights_array(71) := "1100110001";
      weights_array(72) := "1001011101";
      weights_array(73) := "1010000010";
      weights_array(74) := "1101000101";
      weights_array(75) := "0100111011";
      weights_array(76) := "0010110111";
      weights_array(77) := "1000001111";
      weights_array(78) := "0011101010";
      weights_array(79) := "1001110101";
      weights_array(80) := "1110001110";
      weights_array(81) := "0011100110";
      weights_array(82) := "1000111010";
      weights_array(83) := "1000111100";
      weights_array(84) := "1010011001";
      weights_array(85) := "0111100001";
      weights_array(86) := "0101010101";
      weights_array(87) := "1011110100";
      weights_array(88) := "0000011100";
      weights_array(89) := "0001000101";
      weights_array(90) := "1011000100";
      weights_array(91) := "1001001111";
      weights_array(92) := "1010101001";
      weights_array(93) := "0010100101";
      weights_array(94) := "0001001111";
      weights_array(95) := "1001101011";
      weights_array(96) := "1111100101";
      weights_array(97) := "1011100100";
      weights_array(98) := "1010100100";
      weights_array(99) := "0111110100";
      weights_array(100) := "0110000111";
      weights_array(101) := "1010000100";
      weights_array(102) := "0011001100";
      weights_array(103) := "1110100011";
      weights_array(104) := "0100110101";
      weights_array(105) := "0001010011";
      weights_array(106) := "0011000101";
      weights_array(107) := "1111000001";
      weights_array(108) := "1011011011";
      weights_array(109) := "1000101011";
      weights_array(110) := "0111110010";
      weights_array(111) := "1111000101";
      weights_array(112) := "0101110001";
      weights_array(113) := "1010101011";
      weights_array(114) := "0011011000";
      weights_array(115) := "1110111001";
      weights_array(116) := "0100001111";
      weights_array(117) := "0000010010";
      weights_array(118) := "0011010001";
      weights_array(119) := "1010011010";
      weights_array(120) := "1010101011";
      weights_array(121) := "1111010100";
      weights_array(122) := "0110011100";
      weights_array(123) := "0101011010";
      weights_array(124) := "1100110101";
      weights_array(125) := "1011011000";
      weights_array(126) := "1101001101";
      weights_array(127) := "0101100100";
      weights_array(128) := "0110010110";
      weights_array(129) := "1110101100";
      weights_array(130) := "1011000110";
      weights_array(131) := "0000100110";
      weights_array(132) := "0010100000";
      weights_array(133) := "0101010010";
      weights_array(134) := "1001011010";
      weights_array(135) := "0010101010";
      weights_array(136) := "0001111011";
      weights_array(137) := "0101011000";
      weights_array(138) := "1010000111";
      weights_array(139) := "1110011100";
      weights_array(140) := "1000101011";
      weights_array(141) := "0110110111";
      weights_array(142) := "1011010110";
      weights_array(143) := "1001100110";
      weights_array(144) := "0001101011";
      weights_array(145) := "1000100111";
      weights_array(146) := "0101101001";
      weights_array(147) := "0001100011";
      weights_array(148) := "1110101100";
      weights_array(149) := "0000110011";
      weights_array(150) := "0001111011";
      weights_array(151) := "0011100100";
      weights_array(152) := "0011001011";
      weights_array(153) := "1001010110";
      weights_array(154) := "1110110010";
      weights_array(155) := "0101100011";
      weights_array(156) := "0110101000";
      weights_array(157) := "0001110011";
      weights_array(158) := "1110001010";
      weights_array(159) := "0100101100";
      weights_array(160) := "0101010000";
      weights_array(161) := "0111001110";
      weights_array(162) := "0011010101";
      weights_array(163) := "1110010110";
      weights_array(164) := "0011001110";
      weights_array(165) := "0100011101";
      weights_array(166) := "1100011001";
      weights_array(167) := "1010001101";
      weights_array(168) := "0110001100";
      weights_array(169) := "0110110011";
      weights_array(170) := "1001010111";
      weights_array(171) := "0101100100";
      weights_array(172) := "0101100110";
      weights_array(173) := "0001000011";
      weights_array(174) := "0101100011";
      weights_array(175) := "0001111011";
      weights_array(176) := "0010101100";
      weights_array(177) := "1010000100";
      weights_array(178) := "0000111011";
      weights_array(179) := "0110011000";
      weights_array(180) := "0001110010";
      weights_array(181) := "1100011011";
      weights_array(182) := "0110101011";
      weights_array(183) := "0000111010";
      weights_array(184) := "0010111100";
      weights_array(185) := "0101100111";
      weights_array(186) := "0010100110";
      weights_array(187) := "1100111011";
      weights_array(188) := "0011000110";
      weights_array(189) := "1110001001";
      weights_array(190) := "0110001110";
      weights_array(191) := "1010110011";
      weights_array(192) := "1110100001";
      weights_array(193) := "0010110010";
      weights_array(194) := "0010010010";
      weights_array(195) := "1011001001";
      weights_array(196) := "0111101011";
      weights_array(197) := "0111100110";
      weights_array(198) := "0111100010";
      weights_array(199) := "1001011000";
      weights_array(200) := "0000110001";
      weights_array(201) := "1111000100";
      weights_array(202) := "0100101110";
      weights_array(203) := "0111000010";
      weights_array(204) := "0110101011";
      weights_array(205) := "1100000001";
      weights_array(206) := "0111101100";
      weights_array(207) := "0010010110";
      weights_array(208) := "1110110010";
      weights_array(209) := "0010110010";
      weights_array(210) := "1001010111";
      weights_array(211) := "0110101110";
      weights_array(212) := "0010101010";
      weights_array(213) := "0001011010";
      weights_array(214) := "1001000111";
      weights_array(215) := "0110010001";
      weights_array(216) := "1001101100";
      weights_array(217) := "0110000010";
      weights_array(218) := "0010110010";
      weights_array(219) := "0000001111";
      weights_array(220) := "0110101110";
      weights_array(221) := "1100011100";
      weights_array(222) := "1011100001";
      weights_array(223) := "0010110100";
      weights_array(224) := "0010101000";
      weights_array(225) := "0010100110";
      weights_array(226) := "0101010101";
      weights_array(227) := "1110000100";
      weights_array(228) := "1010110010";
      weights_array(229) := "0010001010";
      weights_array(230) := "1001011111";
      weights_array(231) := "0111011110";
      weights_array(232) := "1110010001";
      weights_array(233) := "0101111001";
      weights_array(234) := "0000110011";
      weights_array(235) := "0001001011";
      weights_array(236) := "0010110101";
      weights_array(237) := "1111100000";
      weights_array(238) := "1100100101";
      weights_array(239) := "0100011011";
      weights_array(240) := "0010111010";
      weights_array(241) := "1010011010";
      weights_array(242) := "1110100011";
      weights_array(243) := "1001100101";
      weights_array(244) := "0101101100";
      weights_array(245) := "0010101101";
      weights_array(246) := "1001111011";
      weights_array(247) := "0010100101";
      weights_array(248) := "0011110000";
      weights_array(249) := "0000111001";
      weights_array(250) := "0000110110";
      weights_array(251) := "0010111111";
      weights_array(252) := "1100111011";
      weights_array(253) := "1100001101";
      weights_array(254) := "1000100111";
      weights_array(255) := "1010011100";
      weights_array(256) := "0100110010";
      weights_array(257) := "0101100111";
      weights_array(258) := "1011111100";
      weights_array(259) := "0001110101";
      weights_array(260) := "1000101100";
      weights_array(261) := "0011010111";
      weights_array(262) := "0101101010";
      weights_array(263) := "0000110010";
      weights_array(264) := "0100011011";
      weights_array(265) := "1100011001";
      weights_array(266) := "1100101011";
      weights_array(267) := "1000101110";
      weights_array(268) := "1001001111";
      weights_array(269) := "1001101000";
      weights_array(270) := "1111000111";
      weights_array(271) := "1000100111";
      weights_array(272) := "1100011011";
      weights_array(273) := "0110110001";
      weights_array(274) := "0001100111";
      weights_array(275) := "0111110011";
      weights_array(276) := "1000011011";
      weights_array(277) := "0101100100";
      weights_array(278) := "0011010010";
      weights_array(279) := "0110111001";
      weights_array(280) := "0110100101";
      weights_array(281) := "1110100101";
      weights_array(282) := "0011101110";
      weights_array(283) := "0110011000";
      weights_array(284) := "1000100100";
      weights_array(285) := "0100010101";
      weights_array(286) := "0011011101";
      weights_array(287) := "1110011101";
      weights_array(288) := "0010010010";
      weights_array(289) := "1011000011";
      weights_array(290) := "1111010001";
      weights_array(291) := "0101011001";
      weights_array(292) := "1010011000";
      weights_array(293) := "0100101011";
      weights_array(294) := "1011011010";
      weights_array(295) := "1010101101";
      weights_array(296) := "0111100101";
      weights_array(297) := "1101000011";
      weights_array(298) := "1100100100";
      weights_array(299) := "1010101110";
      weights_array(300) := "0000000000";
      weights_array(301) := "1010010110";
      weights_array(302) := "1011010101";
      weights_array(303) := "0001111100";
      weights_array(304) := "1100001011";
      weights_array(305) := "0101111110";
      weights_array(306) := "0011101000";
      weights_array(307) := "0010000111";
      weights_array(308) := "0101111100";
      weights_array(309) := "0011100001";
      weights_array(310) := "1001100110";
      weights_array(311) := "0011100011";
      weights_array(312) := "1011000111";
      weights_array(313) := "1011001110";
      weights_array(314) := "0111100100";
      weights_array(315) := "0101001011";
      weights_array(316) := "1111111100";
      weights_array(317) := "0000100110";
      weights_array(318) := "0110001000";
      weights_array(319) := "0000101011";
      weights_array(320) := "0101001111";
      weights_array(321) := "0001110100";
      weights_array(322) := "0001111100";
      weights_array(323) := "0111000111";
      weights_array(324) := "1010011011";
      weights_array(325) := "0010011110";
      weights_array(326) := "1111000000";
      weights_array(327) := "0100100110";
      weights_array(328) := "0101011110";
      weights_array(329) := "1000100110";
      weights_array(330) := "1110101000";
      weights_array(331) := "0111010010";
      weights_array(332) := "1101010111";
      weights_array(333) := "1010001111";
      weights_array(334) := "1011100011";
      weights_array(335) := "0000011000";
      weights_array(336) := "0101100110";
      weights_array(337) := "1010101100";
      weights_array(338) := "0101110111";
      weights_array(339) := "1000011100";
      weights_array(340) := "0101111000";
      weights_array(341) := "1100101001";
      weights_array(342) := "1011001011";
      weights_array(343) := "1100101000";
      weights_array(344) := "0110001100";
      weights_array(345) := "0010100111";
      weights_array(346) := "1100101010";
      weights_array(347) := "1111000000";
      weights_array(348) := "1010011111";
      weights_array(349) := "0011001011";
      weights_array(350) := "0100110110";
      weights_array(351) := "1100101010";
      weights_array(352) := "0100101011";
      weights_array(353) := "1111000000";
      weights_array(354) := "0001101100";
      weights_array(355) := "1001000011";
      weights_array(356) := "0100010100";
      weights_array(357) := "0001101101";
      weights_array(358) := "1110011010";
      weights_array(359) := "1010110010";
      weights_array(360) := "0011010011";
      weights_array(361) := "0000110101";
      weights_array(362) := "1110110100";
      weights_array(363) := "0110100011";
      weights_array(364) := "1001110111";
      weights_array(365) := "1110001110";
      weights_array(366) := "0101110101";
      weights_array(367) := "1001000010";
      weights_array(368) := "1010101001";
      weights_array(369) := "0011000101";
      weights_array(370) := "0101110100";
      weights_array(371) := "0000000011";
      weights_array(372) := "0111100100";
      weights_array(373) := "1011110010";
      weights_array(374) := "1010011100";
      weights_array(375) := "0111000011";
      weights_array(376) := "0110100110";
      weights_array(377) := "1101110101";
      weights_array(378) := "0001110011";
      weights_array(379) := "1110010001";
      weights_array(380) := "1011000000";
      weights_array(381) := "0010101110";
      weights_array(382) := "1001011010";
      weights_array(383) := "0001100101";
      weights_array(384) := "1101011111";
      weights_array(385) := "1111100100";
      weights_array(386) := "0001000101";
      weights_array(387) := "1010110010";
      weights_array(388) := "1001111111";
      weights_array(389) := "1101000011";
      weights_array(390) := "0001111001";
      weights_array(391) := "0110100000";
      weights_array(392) := "1000011010";
      weights_array(393) := "0100011011";
      weights_array(394) := "0101010010";
      weights_array(395) := "1010010011";
      weights_array(396) := "1111010010";
      weights_array(397) := "1111010000";
      weights_array(398) := "0011101010";
      weights_array(399) := "0001011100";
      weights_array(400) := "0010100000";
      weights_array(401) := "1111011101";
      weights_array(402) := "0010010010";
      weights_array(403) := "0001011001";
      weights_array(404) := "1011101101";
      weights_array(405) := "0101010101";
      weights_array(406) := "0110000110";
      weights_array(407) := "1000111010";
      weights_array(408) := "1101110011";
      weights_array(409) := "1111000101";
      weights_array(410) := "0111101111";
      weights_array(411) := "1101100101";
      weights_array(412) := "1100011001";
      weights_array(413) := "1011000011";
      weights_array(414) := "0110110001";
      weights_array(415) := "0101100111";
      weights_array(416) := "0010101010";
      weights_array(417) := "1010000101";
      weights_array(418) := "1110000010";
      weights_array(419) := "0111001110";
      weights_array(420) := "0001101110";
      weights_array(421) := "1010011000";
      weights_array(422) := "0001000011";
      weights_array(423) := "1100011001";
      weights_array(424) := "0101011010";
      weights_array(425) := "0100000011";
      weights_array(426) := "0111100001";
      weights_array(427) := "1011000011";
      weights_array(428) := "1001011101";
      weights_array(429) := "1010001101";
      weights_array(430) := "1011001011";
      weights_array(431) := "0111001011";
      weights_array(432) := "0001000110";
      weights_array(433) := "1001010011";
      weights_array(434) := "0110101100";
      weights_array(435) := "1001110001";
      weights_array(436) := "0001010011";
      weights_array(437) := "1010101000";
      weights_array(438) := "1100111010";
      weights_array(439) := "0111011000";
      weights_array(440) := "0000101001";
      weights_array(441) := "0101111000";
      weights_array(442) := "1001011101";
      weights_array(443) := "0010110111";
      weights_array(444) := "1110100101";
      weights_array(445) := "1000101001";
      weights_array(446) := "0000100110";
      weights_array(447) := "1101011100";
      weights_array(448) := "1101001011";
      weights_array(449) := "0000011110";
      weights_array(450) := "0000000111";
      weights_array(451) := "1100011010";
      weights_array(452) := "0001010111";
      weights_array(453) := "0110110101";
      weights_array(454) := "0000011011";
      weights_array(455) := "1100001011";
      weights_array(456) := "1000101011";
      weights_array(457) := "0100100101";
      weights_array(458) := "0101100100";
      weights_array(459) := "1111100011";
      weights_array(460) := "0100111001";
      weights_array(461) := "1100110100";
      weights_array(462) := "1000101110";
      weights_array(463) := "0100011011";
      weights_array(464) := "1010110100";
      weights_array(465) := "0101000010";
      weights_array(466) := "1001000110";
      weights_array(467) := "1000010101";
      weights_array(468) := "0111001001";
      weights_array(469) := "1111000101";
      weights_array(470) := "0110011100";
      weights_array(471) := "0111100011";
      weights_array(472) := "1110101100";
      weights_array(473) := "1011011101";
      weights_array(474) := "1110100110";
      weights_array(475) := "1110001111";
      weights_array(476) := "1000111110";
      weights_array(477) := "0101100010";
      weights_array(478) := "0111100100";
      weights_array(479) := "0011110001";
      weights_array(480) := "0001001110";
      weights_array(481) := "1010001110";
      weights_array(482) := "0100001011";
      weights_array(483) := "0011110001";
      weights_array(484) := "0111001100";
      weights_array(485) := "1000111010";
      weights_array(486) := "0111111000";
      weights_array(487) := "0010110110";
      weights_array(488) := "1010011101";
      weights_array(489) := "0111110000";
      weights_array(490) := "0100111010";
      weights_array(491) := "1100010100";
      weights_array(492) := "1111000101";
      weights_array(493) := "1101000101";
      weights_array(494) := "0100100111";
      weights_array(495) := "0101011100";
      weights_array(496) := "1011101000";
      weights_array(497) := "1001010100";
      weights_array(498) := "0110000011";
      weights_array(499) := "1001011101";
      weights_array(500) := "1000011001";
      weights_array(501) := "1000011011";
      weights_array(502) := "0011101100";
      weights_array(503) := "1010110111";
      weights_array(504) := "1010101001";
      weights_array(505) := "0110011100";
      weights_array(506) := "1100000101";
      weights_array(507) := "0010111100";
      weights_array(508) := "0111011010";
      weights_array(509) := "0101011000";
      weights_array(510) := "0100001011";
      weights_array(511) := "1011101001";
      weights_array(512) := "0000111000";
      weights_array(513) := "0001110011";
      weights_array(514) := "0001100010";
      weights_array(515) := "0011110110";
      weights_array(516) := "1100111011";
      weights_array(517) := "1110100010";
      weights_array(518) := "0110111100";
      weights_array(519) := "0001100011";
      weights_array(520) := "1110000011";
      weights_array(521) := "0111010100";
      weights_array(522) := "0001110011";
      weights_array(523) := "1010001110";
      weights_array(524) := "1001100110";
      weights_array(525) := "1100000111";
      weights_array(526) := "0111010101";
      weights_array(527) := "1110100100";
      weights_array(528) := "0001111101";
      weights_array(529) := "0101110001";
      weights_array(530) := "1100001100";
      weights_array(531) := "1101101001";
      weights_array(532) := "1000011110";
      weights_array(533) := "1001110001";
      weights_array(534) := "1000011010";
      weights_array(535) := "0110000000";
      weights_array(536) := "1000010011";
      weights_array(537) := "1000010111";
      weights_array(538) := "1000011100";
      weights_array(539) := "0011110100";
      weights_array(540) := "0010010011";
      weights_array(541) := "0011000101";
      weights_array(542) := "0001110000";
      weights_array(543) := "0001000101";
      weights_array(544) := "1100101101";
      weights_array(545) := "0100101000";
      weights_array(546) := "0000011011";
      weights_array(547) := "0111000101";
      weights_array(548) := "0110100100";
      weights_array(549) := "0111010010";
      weights_array(550) := "0001001001";
      weights_array(551) := "1100111010";
      weights_array(552) := "1000101111";
      weights_array(553) := "1100100000";
      weights_array(554) := "1101011010";
      weights_array(555) := "0110011101";
      weights_array(556) := "1101001101";
      weights_array(557) := "1010101011";
      weights_array(558) := "1101101010";
      weights_array(559) := "1001010111";
      weights_array(560) := "0011111000";
      weights_array(561) := "0101000110";
      weights_array(562) := "1100000011";
      weights_array(563) := "1101101000";
      weights_array(564) := "0010011111";
      weights_array(565) := "0001000111";
      weights_array(566) := "1111001001";
      weights_array(567) := "0000011011";
      weights_array(568) := "0110100010";
      weights_array(569) := "0111110000";
      weights_array(570) := "1001100101";
      weights_array(571) := "0100111110";
      weights_array(572) := "1000110001";
      weights_array(573) := "1000011010";
      weights_array(574) := "1100100000";
      weights_array(575) := "0111101000";
      weights_array(576) := "0111010101";
      weights_array(577) := "0110100111";
      weights_array(578) := "1000110010";
      weights_array(579) := "0110110010";
      weights_array(580) := "1011100100";
      weights_array(581) := "1100000101";
      weights_array(582) := "1010100011";
      weights_array(583) := "0000101011";
      weights_array(584) := "1100110001";
      weights_array(585) := "1000101111";
      weights_array(586) := "1111100001";
      weights_array(587) := "1000101111";
      weights_array(588) := "0111000101";
      weights_array(589) := "0111101010";
      weights_array(590) := "1001001111";
      weights_array(591) := "0001101011";
      weights_array(592) := "0000101010";
      weights_array(593) := "1101010101";
      weights_array(594) := "1000101011";
      weights_array(595) := "0000111100";
      weights_array(596) := "0101111000";
      weights_array(597) := "1010100011";
      weights_array(598) := "1001001010";
      weights_array(599) := "1111001010";
      weights_array(600) := "1001011100";
      weights_array(601) := "1110000111";
      weights_array(602) := "1010111010";
      weights_array(603) := "0000011011";
      weights_array(604) := "1001110110";
      weights_array(605) := "0101010110";
      weights_array(606) := "0010011111";
      weights_array(607) := "1111000000";

      return weights_array;
    end function;
end fc2_weights_package;

