library ieee;

use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.math_real.all;

use std.textio.all;
use ieee.std_logic_textio.all;


package fc2_weights_package is
    constant HIDDEN_SIZE : integer := 1024;
    constant OUTPUT_SIZE : integer := 10;

    type weights_2_type is array(0 to HIDDEN_SIZE - 1) of std_logic_vector(0 to OUTPUT_SIZE - 1);

    function read_and_populate_weights_2 return weights_2_type;
end fc2_weights_package;

package body fc2_weights_package is
    -- populate the weights_1 array
    function read_and_populate_weights_2 return weights_2_type is
      variable weights_array : weights_2_type;

      variable i : integer := 0;
    begin

      -- weights array: 1024 x 768 
      -- weights_array(0) := "....";
            weights_array(0) := "0010111110";
      weights_array(1) := "0111111100";
      weights_array(2) := "0000011010";
      weights_array(3) := "0110010011";
      weights_array(4) := "0101000110";
      weights_array(5) := "1111010100";
      weights_array(6) := "1001010111";
      weights_array(7) := "1001100111";
      weights_array(8) := "1110001100";
      weights_array(9) := "0101010001";
      weights_array(10) := "0110010101";
      weights_array(11) := "0101110011";
      weights_array(12) := "1000000011";
      weights_array(13) := "0001111011";
      weights_array(14) := "1101110110";
      weights_array(15) := "1010101111";
      weights_array(16) := "0100111100";
      weights_array(17) := "1011001101";
      weights_array(18) := "1110110000";
      weights_array(19) := "0011001011";
      weights_array(20) := "0101101011";
      weights_array(21) := "1110101100";
      weights_array(22) := "1010001001";
      weights_array(23) := "0100010011";
      weights_array(24) := "1111010011";
      weights_array(25) := "0100010011";
      weights_array(26) := "0111010010";
      weights_array(27) := "1101000101";
      weights_array(28) := "0110101000";
      weights_array(29) := "0110000101";
      weights_array(30) := "0110011010";
      weights_array(31) := "1111000100";
      weights_array(32) := "0100001110";
      weights_array(33) := "1100100100";
      weights_array(34) := "0101110100";
      weights_array(35) := "1000111000";
      weights_array(36) := "1100111100";
      weights_array(37) := "1000100100";
      weights_array(38) := "0000011010";
      weights_array(39) := "1110100110";
      weights_array(40) := "1010100000";
      weights_array(41) := "1011100011";
      weights_array(42) := "1110001001";
      weights_array(43) := "0010010011";
      weights_array(44) := "1010111100";
      weights_array(45) := "1000011111";
      weights_array(46) := "1100000101";
      weights_array(47) := "0111101000";
      weights_array(48) := "0110100100";
      weights_array(49) := "0110100010";
      weights_array(50) := "0110100100";
      weights_array(51) := "0000111010";
      weights_array(52) := "1010110000";
      weights_array(53) := "0101010011";
      weights_array(54) := "1110110110";
      weights_array(55) := "1000111010";
      weights_array(56) := "0000011110";
      weights_array(57) := "0111000001";
      weights_array(58) := "0110110011";
      weights_array(59) := "1001111100";
      weights_array(60) := "1111010100";
      weights_array(61) := "1011001110";
      weights_array(62) := "1101010001";
      weights_array(63) := "0111110011";
      weights_array(64) := "1100001111";
      weights_array(65) := "0110010000";
      weights_array(66) := "0101100101";
      weights_array(67) := "0101001111";
      weights_array(68) := "1010010110";
      weights_array(69) := "0110111010";
      weights_array(70) := "0110010000";
      weights_array(71) := "0010010101";
      weights_array(72) := "1010111011";
      weights_array(73) := "1010101000";
      weights_array(74) := "0010100111";
      weights_array(75) := "0101011001";
      weights_array(76) := "1000111110";
      weights_array(77) := "0101011000";
      weights_array(78) := "1001101011";
      weights_array(79) := "1100001001";
      weights_array(80) := "0010101101";
      weights_array(81) := "0111011010";
      weights_array(82) := "0111010101";
      weights_array(83) := "1010111110";
      weights_array(84) := "0000011011";
      weights_array(85) := "0010011001";
      weights_array(86) := "1000011011";
      weights_array(87) := "0110010001";
      weights_array(88) := "0001011100";
      weights_array(89) := "1011000101";
      weights_array(90) := "0001111100";
      weights_array(91) := "0011010000";
      weights_array(92) := "1111110000";
      weights_array(93) := "1100000011";
      weights_array(94) := "1110001011";
      weights_array(95) := "1100011001";
      weights_array(96) := "0100101001";
      weights_array(97) := "0101000111";
      weights_array(98) := "0000110110";
      weights_array(99) := "0001110101";
      weights_array(100) := "0010011011";
      weights_array(101) := "1101111101";
      weights_array(102) := "0110010011";
      weights_array(103) := "1110011100";
      weights_array(104) := "1101101010";
      weights_array(105) := "1110011001";
      weights_array(106) := "1100101100";
      weights_array(107) := "0101110101";
      weights_array(108) := "0011111100";
      weights_array(109) := "1111011001";
      weights_array(110) := "0111100100";
      weights_array(111) := "0001011100";
      weights_array(112) := "1000100001";
      weights_array(113) := "0011001000";
      weights_array(114) := "1110101100";
      weights_array(115) := "0111010101";
      weights_array(116) := "1110100100";
      weights_array(117) := "1001011010";
      weights_array(118) := "0010001111";
      weights_array(119) := "0011100100";
      weights_array(120) := "0100100011";
      weights_array(121) := "0110111110";
      weights_array(122) := "0101110111";
      weights_array(123) := "1101001011";
      weights_array(124) := "0110101111";
      weights_array(125) := "1011100100";
      weights_array(126) := "0010001011";
      weights_array(127) := "0111000010";
      weights_array(128) := "0001010111";
      weights_array(129) := "1100010100";
      weights_array(130) := "1101010101";
      weights_array(131) := "0000010110";
      weights_array(132) := "1010001101";
      weights_array(133) := "1101111001";
      weights_array(134) := "0110011000";
      weights_array(135) := "0101101000";
      weights_array(136) := "0000101110";
      weights_array(137) := "0010010111";
      weights_array(138) := "1000101100";
      weights_array(139) := "0100100011";
      weights_array(140) := "0001100011";
      weights_array(141) := "0100111010";
      weights_array(142) := "1010111111";
      weights_array(143) := "1000110110";
      weights_array(144) := "1100101010";
      weights_array(145) := "0110010011";
      weights_array(146) := "1100011000";
      weights_array(147) := "1000100101";
      weights_array(148) := "1110001100";
      weights_array(149) := "0011110011";
      weights_array(150) := "0011110101";
      weights_array(151) := "1110001110";
      weights_array(152) := "0100100100";
      weights_array(153) := "0101010110";
      weights_array(154) := "1110000011";
      weights_array(155) := "1011100011";
      weights_array(156) := "1000110111";
      weights_array(157) := "0000011011";
      weights_array(158) := "0111011011";
      weights_array(159) := "1001011110";
      weights_array(160) := "1001111010";
      weights_array(161) := "0101110101";
      weights_array(162) := "1111100010";
      weights_array(163) := "1111100111";
      weights_array(164) := "0000011011";
      weights_array(165) := "1000100110";
      weights_array(166) := "1011011101";
      weights_array(167) := "0111011001";
      weights_array(168) := "1001011011";
      weights_array(169) := "0011100001";
      weights_array(170) := "0101100111";
      weights_array(171) := "0101000101";
      weights_array(172) := "1001111001";
      weights_array(173) := "0000101110";
      weights_array(174) := "0101111001";
      weights_array(175) := "0011101001";
      weights_array(176) := "1010010001";
      weights_array(177) := "1100110011";
      weights_array(178) := "1110011101";
      weights_array(179) := "1011100010";
      weights_array(180) := "1000111010";
      weights_array(181) := "0111110110";
      weights_array(182) := "1001011111";
      weights_array(183) := "0110010001";
      weights_array(184) := "0111010110";
      weights_array(185) := "0110011001";
      weights_array(186) := "1010011100";
      weights_array(187) := "1110111010";
      weights_array(188) := "1101001000";
      weights_array(189) := "1001111101";
      weights_array(190) := "0101010010";
      weights_array(191) := "1001001111";
      weights_array(192) := "0101100100";
      weights_array(193) := "0000110010";
      weights_array(194) := "1100001001";
      weights_array(195) := "0110001011";
      weights_array(196) := "1010001100";
      weights_array(197) := "0001110011";
      weights_array(198) := "1001110001";
      weights_array(199) := "0011111000";
      weights_array(200) := "1011110001";
      weights_array(201) := "0001100011";
      weights_array(202) := "1011000101";
      weights_array(203) := "0101011100";
      weights_array(204) := "1000011011";
      weights_array(205) := "0110001010";
      weights_array(206) := "0111000110";
      weights_array(207) := "0011110000";
      weights_array(208) := "1000011011";
      weights_array(209) := "0000111101";
      weights_array(210) := "0011010010";
      weights_array(211) := "1010110001";
      weights_array(212) := "0010010110";
      weights_array(213) := "1100101010";
      weights_array(214) := "1111101001";
      weights_array(215) := "0111011000";
      weights_array(216) := "1110100001";
      weights_array(217) := "0100101110";
      weights_array(218) := "0110101000";
      weights_array(219) := "1011100110";
      weights_array(220) := "1001010111";
      weights_array(221) := "1100100100";
      weights_array(222) := "1111100100";
      weights_array(223) := "1100110001";
      weights_array(224) := "0001001011";
      weights_array(225) := "1110010000";
      weights_array(226) := "1101010110";
      weights_array(227) := "0110010111";
      weights_array(228) := "1101010110";
      weights_array(229) := "1110011000";
      weights_array(230) := "0111001001";
      weights_array(231) := "0101100110";
      weights_array(232) := "1110000011";
      weights_array(233) := "0011000100";
      weights_array(234) := "1000101011";
      weights_array(235) := "0001011101";
      weights_array(236) := "0010010001";
      weights_array(237) := "1010101001";
      weights_array(238) := "0011001110";
      weights_array(239) := "1101101110";
      weights_array(240) := "1110000111";
      weights_array(241) := "0100110011";
      weights_array(242) := "0101110100";
      weights_array(243) := "1111110100";
      weights_array(244) := "1010011010";
      weights_array(245) := "0010011101";
      weights_array(246) := "0111001001";
      weights_array(247) := "1010010101";
      weights_array(248) := "1000100111";
      weights_array(249) := "1100010111";
      weights_array(250) := "1111000011";
      weights_array(251) := "1010001101";
      weights_array(252) := "0111100010";
      weights_array(253) := "1001010101";
      weights_array(254) := "1111000100";
      weights_array(255) := "0110111101";
      weights_array(256) := "0011010000";
      weights_array(257) := "0110101110";
      weights_array(258) := "0001000011";
      weights_array(259) := "1111010011";
      weights_array(260) := "1001111100";
      weights_array(261) := "1011010101";
      weights_array(262) := "1110010100";
      weights_array(263) := "1001001011";
      weights_array(264) := "1001100111";
      weights_array(265) := "1101110100";
      weights_array(266) := "1000001011";
      weights_array(267) := "0001110100";
      weights_array(268) := "1100001100";
      weights_array(269) := "0110010011";
      weights_array(270) := "0010101110";
      weights_array(271) := "0101000111";
      weights_array(272) := "0000110110";
      weights_array(273) := "0111011100";
      weights_array(274) := "0111011010";
      weights_array(275) := "0110110100";
      weights_array(276) := "1010110001";
      weights_array(277) := "0000101100";
      weights_array(278) := "1110111010";
      weights_array(279) := "0011111000";
      weights_array(280) := "1110001011";
      weights_array(281) := "0100110111";
      weights_array(282) := "0011010000";
      weights_array(283) := "1111010000";
      weights_array(284) := "1010100111";
      weights_array(285) := "0110010000";
      weights_array(286) := "1010101010";
      weights_array(287) := "0111111111";
      weights_array(288) := "0110100011";
      weights_array(289) := "0001100110";
      weights_array(290) := "0000100001";
      weights_array(291) := "0111101100";
      weights_array(292) := "1000001101";
      weights_array(293) := "0100001000";
      weights_array(294) := "0000101001";
      weights_array(295) := "0010011010";
      weights_array(296) := "1001010100";
      weights_array(297) := "0001100001";
      weights_array(298) := "0011000110";
      weights_array(299) := "1000001110";
      weights_array(300) := "1110000101";
      weights_array(301) := "0000110111";
      weights_array(302) := "1000010110";
      weights_array(303) := "1011100100";
      weights_array(304) := "0111100001";
      weights_array(305) := "1011001001";
      weights_array(306) := "1000100111";
      weights_array(307) := "0011101101";
      weights_array(308) := "0000010101";
      weights_array(309) := "1000111110";
      weights_array(310) := "0100001001";
      weights_array(311) := "1110000001";
      weights_array(312) := "1000110101";
      weights_array(313) := "0111000010";
      weights_array(314) := "1111001111";
      weights_array(315) := "1101100110";
      weights_array(316) := "1011101101";
      weights_array(317) := "1111100011";
      weights_array(318) := "0101110100";
      weights_array(319) := "0110011100";
      weights_array(320) := "0011111110";
      weights_array(321) := "1111000110";
      weights_array(322) := "0011010110";
      weights_array(323) := "1010001100";
      weights_array(324) := "1001100101";
      weights_array(325) := "1110001010";
      weights_array(326) := "1110100111";
      weights_array(327) := "0110000111";
      weights_array(328) := "1010110010";
      weights_array(329) := "1100110110";
      weights_array(330) := "1100111010";
      weights_array(331) := "0000011011";
      weights_array(332) := "1101010100";
      weights_array(333) := "0011011111";
      weights_array(334) := "1111101000";
      weights_array(335) := "1101010100";
      weights_array(336) := "1101100011";
      weights_array(337) := "1000011110";
      weights_array(338) := "0110011110";
      weights_array(339) := "0010100111";
      weights_array(340) := "0011010100";
      weights_array(341) := "1001001011";
      weights_array(342) := "0001010101";
      weights_array(343) := "0101100111";
      weights_array(344) := "1000011011";
      weights_array(345) := "1101111000";
      weights_array(346) := "1001001011";
      weights_array(347) := "1010001110";
      weights_array(348) := "1001000011";
      weights_array(349) := "0010010010";
      weights_array(350) := "0001111110";
      weights_array(351) := "1011101001";
      weights_array(352) := "1111010010";
      weights_array(353) := "0011010101";
      weights_array(354) := "1001010101";
      weights_array(355) := "0110001110";
      weights_array(356) := "1011111010";
      weights_array(357) := "1111000100";
      weights_array(358) := "0011110000";
      weights_array(359) := "0010111110";
      weights_array(360) := "0101110110";
      weights_array(361) := "0001000101";
      weights_array(362) := "1001110001";
      weights_array(363) := "1000001110";
      weights_array(364) := "0101011000";
      weights_array(365) := "1010110010";
      weights_array(366) := "1001101011";
      weights_array(367) := "1010110011";
      weights_array(368) := "1010111010";
      weights_array(369) := "1110111011";
      weights_array(370) := "0100101010";
      weights_array(371) := "1001000101";
      weights_array(372) := "1111000100";
      weights_array(373) := "1110101110";
      weights_array(374) := "1001000011";
      weights_array(375) := "0100111001";
      weights_array(376) := "1001011001";
      weights_array(377) := "1111000100";
      weights_array(378) := "0011010001";
      weights_array(379) := "1111010000";
      weights_array(380) := "1001011011";
      weights_array(381) := "1111101110";
      weights_array(382) := "1110011010";
      weights_array(383) := "0011101010";
      weights_array(384) := "1101100100";
      weights_array(385) := "1000110101";
      weights_array(386) := "1111000010";
      weights_array(387) := "0011100101";
      weights_array(388) := "0100011101";
      weights_array(389) := "0010101011";
      weights_array(390) := "1001100111";
      weights_array(391) := "0100111000";
      weights_array(392) := "1010000111";
      weights_array(393) := "0111000001";
      weights_array(394) := "0101000010";
      weights_array(395) := "0011010100";
      weights_array(396) := "0011110011";
      weights_array(397) := "0111111100";
      weights_array(398) := "1010011011";
      weights_array(399) := "1010101100";
      weights_array(400) := "1001100101";
      weights_array(401) := "1000111100";
      weights_array(402) := "0101110011";
      weights_array(403) := "0011010010";
      weights_array(404) := "1010100001";
      weights_array(405) := "0100101011";
      weights_array(406) := "1111001001";
      weights_array(407) := "1110101011";
      weights_array(408) := "0011111011";
      weights_array(409) := "1011110101";
      weights_array(410) := "1010001011";
      weights_array(411) := "1101010100";
      weights_array(412) := "0011001100";
      weights_array(413) := "1111001011";
      weights_array(414) := "0101101100";
      weights_array(415) := "0110001101";
      weights_array(416) := "0001111000";
      weights_array(417) := "0000110011";
      weights_array(418) := "0000111010";
      weights_array(419) := "0101101101";
      weights_array(420) := "0010110101";
      weights_array(421) := "1110011001";
      weights_array(422) := "0111110000";
      weights_array(423) := "1100101110";
      weights_array(424) := "0011000110";
      weights_array(425) := "0000111100";
      weights_array(426) := "1110010100";
      weights_array(427) := "0100000011";
      weights_array(428) := "1100111010";
      weights_array(429) := "1111000110";
      weights_array(430) := "1000010110";
      weights_array(431) := "1101001011";
      weights_array(432) := "1000100101";
      weights_array(433) := "0100001011";
      weights_array(434) := "1010110101";
      weights_array(435) := "1011100101";
      weights_array(436) := "0111100010";
      weights_array(437) := "1110001010";
      weights_array(438) := "1001100101";
      weights_array(439) := "1100101000";
      weights_array(440) := "0101111000";
      weights_array(441) := "0100010011";
      weights_array(442) := "0111010101";
      weights_array(443) := "0111010011";
      weights_array(444) := "0001011110";
      weights_array(445) := "1011011111";
      weights_array(446) := "0010110001";
      weights_array(447) := "0111100000";
      weights_array(448) := "0101010111";
      weights_array(449) := "0011011001";
      weights_array(450) := "0100111010";
      weights_array(451) := "1010011001";
      weights_array(452) := "0110100000";
      weights_array(453) := "0111100101";
      weights_array(454) := "0001110010";
      weights_array(455) := "0111100010";
      weights_array(456) := "0011110101";
      weights_array(457) := "1010011000";
      weights_array(458) := "0111001110";
      weights_array(459) := "1101100001";
      weights_array(460) := "0101100011";
      weights_array(461) := "1011000010";
      weights_array(462) := "0101110011";
      weights_array(463) := "0000011011";
      weights_array(464) := "1011101101";
      weights_array(465) := "0101101010";
      weights_array(466) := "0100010010";
      weights_array(467) := "1111011000";
      weights_array(468) := "1001100011";
      weights_array(469) := "0111001010";
      weights_array(470) := "0101000101";
      weights_array(471) := "1001010010";
      weights_array(472) := "0110011011";
      weights_array(473) := "1100100001";
      weights_array(474) := "1111001001";
      weights_array(475) := "1111101100";
      weights_array(476) := "0001011001";
      weights_array(477) := "1010100001";
      weights_array(478) := "0010100101";
      weights_array(479) := "0110010111";
      weights_array(480) := "1111010100";
      weights_array(481) := "1011001111";
      weights_array(482) := "1001000110";
      weights_array(483) := "1111110100";
      weights_array(484) := "1001111100";
      weights_array(485) := "1010101100";
      weights_array(486) := "1000100101";
      weights_array(487) := "1001010010";
      weights_array(488) := "1011101000";
      weights_array(489) := "0010011010";
      weights_array(490) := "0111101100";
      weights_array(491) := "0110011001";
      weights_array(492) := "0111100011";
      weights_array(493) := "0001111010";
      weights_array(494) := "1000011001";
      weights_array(495) := "0100001111";
      weights_array(496) := "0001000010";
      weights_array(497) := "1001000101";
      weights_array(498) := "0001100011";
      weights_array(499) := "1100111011";
      weights_array(500) := "1001111110";
      weights_array(501) := "0011001011";
      weights_array(502) := "0010100011";
      weights_array(503) := "1110010001";
      weights_array(504) := "1110101001";
      weights_array(505) := "0110111100";
      weights_array(506) := "1111000110";
      weights_array(507) := "0111100110";
      weights_array(508) := "1000010111";
      weights_array(509) := "0000101010";
      weights_array(510) := "1110101000";
      weights_array(511) := "0010000100";
      weights_array(512) := "1111110010";
      weights_array(513) := "1101101011";
      weights_array(514) := "1001110000";
      weights_array(515) := "1100101011";
      weights_array(516) := "0000111100";
      weights_array(517) := "0001101000";
      weights_array(518) := "1101111011";
      weights_array(519) := "0111110101";
      weights_array(520) := "0000100001";
      weights_array(521) := "1001101011";
      weights_array(522) := "0111011010";
      weights_array(523) := "1011011011";
      weights_array(524) := "0110011101";
      weights_array(525) := "0001010110";
      weights_array(526) := "0010001010";
      weights_array(527) := "1100100101";
      weights_array(528) := "1010010001";
      weights_array(529) := "0101011111";
      weights_array(530) := "1111000001";
      weights_array(531) := "0111000000";
      weights_array(532) := "0100111011";
      weights_array(533) := "1001010000";
      weights_array(534) := "1110101111";
      weights_array(535) := "0010111000";
      weights_array(536) := "0111001010";
      weights_array(537) := "0101011100";
      weights_array(538) := "1001100110";
      weights_array(539) := "1111101100";
      weights_array(540) := "1011100101";
      weights_array(541) := "1000000001";
      weights_array(542) := "1011001000";
      weights_array(543) := "0000101011";
      weights_array(544) := "0001100001";
      weights_array(545) := "1010000111";
      weights_array(546) := "1100001101";
      weights_array(547) := "1000010001";
      weights_array(548) := "1111100010";
      weights_array(549) := "1011000100";
      weights_array(550) := "1000110010";
      weights_array(551) := "1101010001";
      weights_array(552) := "0101110100";
      weights_array(553) := "1110011001";
      weights_array(554) := "1100101111";
      weights_array(555) := "1110001001";
      weights_array(556) := "0110000110";
      weights_array(557) := "1001110101";
      weights_array(558) := "1010010111";
      weights_array(559) := "1010001110";
      weights_array(560) := "0101110101";
      weights_array(561) := "0011001100";
      weights_array(562) := "1110100101";
      weights_array(563) := "0011110110";
      weights_array(564) := "1011001100";
      weights_array(565) := "0001000111";
      weights_array(566) := "0100111011";
      weights_array(567) := "0101000110";
      weights_array(568) := "0111000100";
      weights_array(569) := "0010100110";
      weights_array(570) := "1100010010";
      weights_array(571) := "0011100101";
      weights_array(572) := "1011100100";
      weights_array(573) := "1100100101";
      weights_array(574) := "1010101000";
      weights_array(575) := "0111010010";
      weights_array(576) := "0000011011";
      weights_array(577) := "0000101001";
      weights_array(578) := "0111010110";
      weights_array(579) := "0111010100";
      weights_array(580) := "0111010010";
      weights_array(581) := "1011000110";
      weights_array(582) := "0110100111";
      weights_array(583) := "1011001100";
      weights_array(584) := "0101100011";
      weights_array(585) := "0000101110";
      weights_array(586) := "1010100101";
      weights_array(587) := "1101101001";
      weights_array(588) := "0111000011";
      weights_array(589) := "1001100011";
      weights_array(590) := "0001110100";
      weights_array(591) := "1111000101";
      weights_array(592) := "1111100100";
      weights_array(593) := "0101011110";
      weights_array(594) := "0111110110";
      weights_array(595) := "0001111011";
      weights_array(596) := "0110100111";
      weights_array(597) := "0011000110";
      weights_array(598) := "0000110111";
      weights_array(599) := "1011010111";
      weights_array(600) := "1011100011";
      weights_array(601) := "0010111011";
      weights_array(602) := "1111000101";
      weights_array(603) := "1010011110";
      weights_array(604) := "1110111000";
      weights_array(605) := "0100111010";
      weights_array(606) := "0100100011";
      weights_array(607) := "0110011011";
      weights_array(608) := "0110011000";
      weights_array(609) := "0000100111";
      weights_array(610) := "1001100101";
      weights_array(611) := "0111001101";
      weights_array(612) := "1011010111";
      weights_array(613) := "0100101001";
      weights_array(614) := "0011110111";
      weights_array(615) := "1010000110";
      weights_array(616) := "0111101000";
      weights_array(617) := "0100010101";
      weights_array(618) := "0110000011";
      weights_array(619) := "1011101000";
      weights_array(620) := "1100011100";
      weights_array(621) := "1000110010";
      weights_array(622) := "1100111000";
      weights_array(623) := "1000101011";
      weights_array(624) := "0000111110";
      weights_array(625) := "1011111000";
      weights_array(626) := "0001001011";
      weights_array(627) := "1001100110";
      weights_array(628) := "1000110001";
      weights_array(629) := "0100111010";
      weights_array(630) := "1110011101";
      weights_array(631) := "0011011100";
      weights_array(632) := "1001100001";
      weights_array(633) := "0100111110";
      weights_array(634) := "1010100100";
      weights_array(635) := "1011000100";
      weights_array(636) := "1111010010";
      weights_array(637) := "1100110111";
      weights_array(638) := "0011100101";
      weights_array(639) := "1010011100";
      weights_array(640) := "0101101100";
      weights_array(641) := "1011001010";
      weights_array(642) := "1111001001";
      weights_array(643) := "0111100100";
      weights_array(644) := "0100110111";
      weights_array(645) := "1110101000";
      weights_array(646) := "0010001100";
      weights_array(647) := "1010001111";
      weights_array(648) := "0111000010";
      weights_array(649) := "0110100001";
      weights_array(650) := "1011100101";
      weights_array(651) := "0001010110";
      weights_array(652) := "1110111000";
      weights_array(653) := "0011101001";
      weights_array(654) := "1101011010";
      weights_array(655) := "1000100110";
      weights_array(656) := "1000101011";
      weights_array(657) := "1111000001";
      weights_array(658) := "1110101101";
      weights_array(659) := "1110010000";
      weights_array(660) := "1101011011";
      weights_array(661) := "1000011101";
      weights_array(662) := "0010100101";
      weights_array(663) := "1101101100";
      weights_array(664) := "0001110100";
      weights_array(665) := "0100101001";
      weights_array(666) := "0110111101";
      weights_array(667) := "0100110100";
      weights_array(668) := "0001101011";
      weights_array(669) := "1001101001";
      weights_array(670) := "1011111001";
      weights_array(671) := "0001100111";
      weights_array(672) := "0111001100";
      weights_array(673) := "0101110011";
      weights_array(674) := "0010011101";
      weights_array(675) := "1001000011";
      weights_array(676) := "0111100000";
      weights_array(677) := "1000111011";
      weights_array(678) := "0101111101";
      weights_array(679) := "1001100100";
      weights_array(680) := "1111000001";
      weights_array(681) := "1001110011";
      weights_array(682) := "0010011111";
      weights_array(683) := "1101110001";
      weights_array(684) := "0100001101";
      weights_array(685) := "0101110100";
      weights_array(686) := "1101000010";
      weights_array(687) := "0110100101";
      weights_array(688) := "1011111100";
      weights_array(689) := "0011111000";
      weights_array(690) := "0110000100";
      weights_array(691) := "0001011010";
      weights_array(692) := "1100111011";
      weights_array(693) := "0001001010";
      weights_array(694) := "0010100110";
      weights_array(695) := "0101011001";
      weights_array(696) := "1110001101";
      weights_array(697) := "0111000011";
      weights_array(698) := "1110001110";
      weights_array(699) := "0100010011";
      weights_array(700) := "0001110111";
      weights_array(701) := "1001101100";
      weights_array(702) := "0111101010";
      weights_array(703) := "0011110010";
      weights_array(704) := "1110101010";
      weights_array(705) := "1111001011";
      weights_array(706) := "1000111000";
      weights_array(707) := "0000101011";
      weights_array(708) := "0101111001";
      weights_array(709) := "0100100011";
      weights_array(710) := "0001110000";
      weights_array(711) := "0000010111";
      weights_array(712) := "1101011110";
      weights_array(713) := "1110000110";
      weights_array(714) := "0001100110";
      weights_array(715) := "0100110000";
      weights_array(716) := "1100011110";
      weights_array(717) := "1110100010";
      weights_array(718) := "1110001100";
      weights_array(719) := "1010111011";
      weights_array(720) := "1010100100";
      weights_array(721) := "1101000111";
      weights_array(722) := "0011010110";
      weights_array(723) := "1101010100";
      weights_array(724) := "0001010011";
      weights_array(725) := "0010101010";
      weights_array(726) := "0000101010";
      weights_array(727) := "0000111011";
      weights_array(728) := "1110100011";
      weights_array(729) := "0101111001";
      weights_array(730) := "1000010001";
      weights_array(731) := "0100101010";
      weights_array(732) := "0100101001";
      weights_array(733) := "1010000001";
      weights_array(734) := "1100110111";
      weights_array(735) := "0101000101";
      weights_array(736) := "1001011011";
      weights_array(737) := "0101101111";
      weights_array(738) := "0100101001";
      weights_array(739) := "1100010100";
      weights_array(740) := "1010001101";
      weights_array(741) := "1010111010";
      weights_array(742) := "0101110111";
      weights_array(743) := "0000110111";
      weights_array(744) := "0000111101";
      weights_array(745) := "0110100100";
      weights_array(746) := "0000100111";
      weights_array(747) := "1010010110";
      weights_array(748) := "0000011001";
      weights_array(749) := "1010110010";
      weights_array(750) := "0011111011";
      weights_array(751) := "1111000110";
      weights_array(752) := "0110100010";
      weights_array(753) := "0000101011";
      weights_array(754) := "1101011010";
      weights_array(755) := "0000000101";
      weights_array(756) := "0101100100";
      weights_array(757) := "1011010100";
      weights_array(758) := "0101011101";
      weights_array(759) := "0001110011";
      weights_array(760) := "0000100110";
      weights_array(761) := "1110000010";
      weights_array(762) := "0011011101";
      weights_array(763) := "0101100011";
      weights_array(764) := "1011011100";
      weights_array(765) := "0001110111";
      weights_array(766) := "0001011010";
      weights_array(767) := "0011000111";
      weights_array(768) := "1000011100";
      weights_array(769) := "1011100000";
      weights_array(770) := "0001010000";
      weights_array(771) := "1011011000";
      weights_array(772) := "0101011010";
      weights_array(773) := "1000100111";
      weights_array(774) := "1101001000";
      weights_array(775) := "1000010100";
      weights_array(776) := "1101001010";
      weights_array(777) := "0001010001";
      weights_array(778) := "0111100011";
      weights_array(779) := "0110111001";
      weights_array(780) := "0101101110";
      weights_array(781) := "1000101101";
      weights_array(782) := "1011010101";
      weights_array(783) := "1010111000";
      weights_array(784) := "1010000110";
      weights_array(785) := "0111010110";
      weights_array(786) := "1010101101";
      weights_array(787) := "1000011010";
      weights_array(788) := "1100001100";
      weights_array(789) := "0111001100";
      weights_array(790) := "1110100001";
      weights_array(791) := "1110101011";
      weights_array(792) := "0101011001";
      weights_array(793) := "1010110010";
      weights_array(794) := "1100001001";
      weights_array(795) := "0101011010";
      weights_array(796) := "1011010001";
      weights_array(797) := "0111011001";
      weights_array(798) := "0010101101";
      weights_array(799) := "1101000001";
      weights_array(800) := "0001010001";
      weights_array(801) := "1100110001";
      weights_array(802) := "1010100110";
      weights_array(803) := "1011001011";
      weights_array(804) := "1010010100";
      weights_array(805) := "1011011101";
      weights_array(806) := "0110110111";
      weights_array(807) := "0101010011";
      weights_array(808) := "0100110010";
      weights_array(809) := "0001010101";
      weights_array(810) := "1001000111";
      weights_array(811) := "0010111011";
      weights_array(812) := "0111001100";
      weights_array(813) := "0001011010";
      weights_array(814) := "0110011001";
      weights_array(815) := "0111000101";
      weights_array(816) := "1101010101";
      weights_array(817) := "0111000110";
      weights_array(818) := "0100110001";
      weights_array(819) := "1000111101";
      weights_array(820) := "1000110110";
      weights_array(821) := "1111010100";
      weights_array(822) := "1100001101";
      weights_array(823) := "1001011000";
      weights_array(824) := "0011101101";
      weights_array(825) := "0101101010";
      weights_array(826) := "0001000110";
      weights_array(827) := "0110010101";
      weights_array(828) := "1100111000";
      weights_array(829) := "0011111001";
      weights_array(830) := "1100100101";
      weights_array(831) := "0110111100";
      weights_array(832) := "1111000110";
      weights_array(833) := "0010001000";
      weights_array(834) := "0110101101";
      weights_array(835) := "1011000101";
      weights_array(836) := "0111010000";
      weights_array(837) := "1001000101";
      weights_array(838) := "0001100001";
      weights_array(839) := "0001111101";
      weights_array(840) := "1001110101";
      weights_array(841) := "1100101011";
      weights_array(842) := "1110110000";
      weights_array(843) := "1000011111";
      weights_array(844) := "1000010100";
      weights_array(845) := "0110011001";
      weights_array(846) := "0100110111";
      weights_array(847) := "0101001001";
      weights_array(848) := "0111000001";
      weights_array(849) := "1111101100";
      weights_array(850) := "1000101011";
      weights_array(851) := "1000101110";
      weights_array(852) := "0110101010";
      weights_array(853) := "0001111000";
      weights_array(854) := "1110101110";
      weights_array(855) := "0010110110";
      weights_array(856) := "1110101011";
      weights_array(857) := "0101111010";
      weights_array(858) := "0000011111";
      weights_array(859) := "1111001011";
      weights_array(860) := "0000101011";
      weights_array(861) := "0110001101";
      weights_array(862) := "0001011011";
      weights_array(863) := "1100011110";
      weights_array(864) := "0010011001";
      weights_array(865) := "1000010000";
      weights_array(866) := "1011011010";
      weights_array(867) := "1001110000";
      weights_array(868) := "0111101011";
      weights_array(869) := "1101010101";
      weights_array(870) := "1011011001";
      weights_array(871) := "0010110011";
      weights_array(872) := "0011110111";
      weights_array(873) := "1010010011";
      weights_array(874) := "1011000110";
      weights_array(875) := "0001111110";
      weights_array(876) := "0001110100";
      weights_array(877) := "1001010111";
      weights_array(878) := "0011011101";
      weights_array(879) := "1010010110";
      weights_array(880) := "1011001010";
      weights_array(881) := "1001010000";
      weights_array(882) := "1111000100";
      weights_array(883) := "0100111001";
      weights_array(884) := "1110101010";
      weights_array(885) := "0001101100";
      weights_array(886) := "1110100000";
      weights_array(887) := "0110001110";
      weights_array(888) := "0100100101";
      weights_array(889) := "0000111111";
      weights_array(890) := "1101010100";
      weights_array(891) := "0100001011";
      weights_array(892) := "0110101010";
      weights_array(893) := "1110101010";
      weights_array(894) := "1101001001";
      weights_array(895) := "0101011100";
      weights_array(896) := "1110100111";
      weights_array(897) := "1101110001";
      weights_array(898) := "0000000111";
      weights_array(899) := "1000001011";
      weights_array(900) := "0111011000";
      weights_array(901) := "0101110101";
      weights_array(902) := "1010111000";
      weights_array(903) := "0001010111";
      weights_array(904) := "1010011001";
      weights_array(905) := "0100111010";
      weights_array(906) := "1101111111";
      weights_array(907) := "0101100100";
      weights_array(908) := "1111101001";
      weights_array(909) := "1011100001";
      weights_array(910) := "0100100110";
      weights_array(911) := "1101100100";
      weights_array(912) := "1111000101";
      weights_array(913) := "0110011100";
      weights_array(914) := "1010010110";
      weights_array(915) := "0100011001";
      weights_array(916) := "0100110001";
      weights_array(917) := "1011011001";
      weights_array(918) := "1010101010";
      weights_array(919) := "0111011010";
      weights_array(920) := "1011111001";
      weights_array(921) := "1000000011";
      weights_array(922) := "0010110001";
      weights_array(923) := "1100001110";
      weights_array(924) := "0111101010";
      weights_array(925) := "1111010101";
      weights_array(926) := "1010111000";
      weights_array(927) := "1001101000";
      weights_array(928) := "0111110110";
      weights_array(929) := "1011101110";
      weights_array(930) := "0111010011";
      weights_array(931) := "1001010010";
      weights_array(932) := "0011111101";
      weights_array(933) := "1010011010";
      weights_array(934) := "0110111100";
      weights_array(935) := "1000011110";
      weights_array(936) := "0101111010";
      weights_array(937) := "0100111010";
      weights_array(938) := "1001101001";
      weights_array(939) := "0111100110";
      weights_array(940) := "1101111110";
      weights_array(941) := "0100010101";
      weights_array(942) := "1011110101";
      weights_array(943) := "0110010111";
      weights_array(944) := "1100101000";
      weights_array(945) := "1101100100";
      weights_array(946) := "1010000011";
      weights_array(947) := "1100011010";
      weights_array(948) := "1111101100";
      weights_array(949) := "1101100110";
      weights_array(950) := "0000011010";
      weights_array(951) := "1110100100";
      weights_array(952) := "1010011110";
      weights_array(953) := "0111100110";
      weights_array(954) := "0110100010";
      weights_array(955) := "0100101110";
      weights_array(956) := "1011101001";
      weights_array(957) := "0011010100";
      weights_array(958) := "1010111000";
      weights_array(959) := "0110011001";
      weights_array(960) := "1111001101";
      weights_array(961) := "0111110010";
      weights_array(962) := "0000101010";
      weights_array(963) := "1100011100";
      weights_array(964) := "0010010001";
      weights_array(965) := "0110110010";
      weights_array(966) := "0110101100";
      weights_array(967) := "0011000011";
      weights_array(968) := "1011100100";
      weights_array(969) := "1001101011";
      weights_array(970) := "0010010010";
      weights_array(971) := "1000111111";
      weights_array(972) := "0001001011";
      weights_array(973) := "1010000101";
      weights_array(974) := "0111010001";
      weights_array(975) := "1010001001";
      weights_array(976) := "1111011100";
      weights_array(977) := "1101100001";
      weights_array(978) := "0101110110";
      weights_array(979) := "0100111010";
      weights_array(980) := "1100011110";
      weights_array(981) := "0101110101";
      weights_array(982) := "1011001101";
      weights_array(983) := "0110011010";
      weights_array(984) := "0101111000";
      weights_array(985) := "0101110011";
      weights_array(986) := "0111100111";
      weights_array(987) := "0001001100";
      weights_array(988) := "1001000100";
      weights_array(989) := "1001100101";
      weights_array(990) := "0011001000";
      weights_array(991) := "1101000110";
      weights_array(992) := "0111010011";
      weights_array(993) := "1001011001";
      weights_array(994) := "1010110001";
      weights_array(995) := "1100101001";
      weights_array(996) := "1010111100";
      weights_array(997) := "1000011001";
      weights_array(998) := "1000101110";
      weights_array(999) := "1100111100";
      weights_array(1000) := "1111001100";
      weights_array(1001) := "0001110111";
      weights_array(1002) := "1110110010";
      weights_array(1003) := "1001010001";
      weights_array(1004) := "1110001110";
      weights_array(1005) := "0001011110";
      weights_array(1006) := "0111000100";
      weights_array(1007) := "1011011000";
      weights_array(1008) := "1001111000";
      weights_array(1009) := "1001010000";
      weights_array(1010) := "0111100001";
      weights_array(1011) := "1110110000";
      weights_array(1012) := "1000011101";
      weights_array(1013) := "0000001110";
      weights_array(1014) := "1110000101";
      weights_array(1015) := "0111001001";
      weights_array(1016) := "0110001010";
      weights_array(1017) := "0111010100";
      weights_array(1018) := "0001001101";
      weights_array(1019) := "0101000111";
      weights_array(1020) := "0110000010";
      weights_array(1021) := "1111110011";
      weights_array(1022) := "1110100000";
      weights_array(1023) := "1111001100";

      return weights_array;
    end function;
end fc2_weights_package;

